module encoder2_1 (
    input wire[1:0] encoder_in;
    output reg[0] encoder_out;
);
    
endmodule